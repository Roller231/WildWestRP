/       D a t a ,   A s s e m b l y - C S h a r p        d a t a G o l d �     d a t a S t o r a g e /      S y s t e m . I n t 3 2 [ ] ,   m s c o r l i b          
   
   d a t a I n c o m e 0                  d a t a M a x I n c o m e 0            
   	   d a t a L e v e l 0                  d a t a U p g r a d e C o s t 0            
      d a t a T i m e E a r n /      S y s t e m . S i n g l e [ ] ,   m s c o r l i b             @   d a t a U p g r a d e G o l d E a r n 0            
      d a t a U p g r a d e N e w M a x I n c o m e 0                  g a m e O b j e c t s /      S y s t e m . S t r i n g [ ] ,   m s c o r l i b 	          (   S c h a h t a ( C l o n e )    p o s X 0   
         PJ�?   p o s Y 0            ��
   i s O c c u p p e d /      S y s t e m . B o o l e a n [ ] ,   m s c o r l i b          	   i n d e x T i l e 0            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              